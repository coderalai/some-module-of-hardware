`include "defines.v"

module clint(
    input   wire            clk,
    input   wire            rst,

    // from core
    input   wire    [`INT_BUS    ]      int_flag_i,

    // from id
    input   wire    [`InstBus     ]      inst_i          ,
    input   wire    [`InstAddrBus]      inst_addr_i     ,

    // from ex
    input   wire                        jump_flag_i     ,
    input   wire    [`InstAddrBus]      jump_addr_i     ,
    input   wire                        div_started_i   ,

    // from ctrl
    input   wire    [`Hold_Flag_Bus]    hold_flag_i     ,

    // from csr_reg
    input   wire    [`RegBus      ]     data_i          ,
    input   wire    [`RegBus      ]     csr_mtvec       ,
    input   wire    [`RegBus      ]     csr_mepc        ,
    input   wire    [`RegBus      ]     csr_mstatus     ,

    input   wire                        global_int_en_i ,

    // to ctrl
    output  wire                        hold_flag_o      ,

    // to csr_reg
    output  reg                         we_o             ,
    output  reg     [`MemAddrBus  ]     waddr_o          ,
    output  reg     [`MemAddrBus  ]     raddr_o          ,
    output  reg     [`RegBus      ]     data_o           ,

    // to ex
    output  reg     [`InstAddrBus]      int_addr_o      ,
    output  reg                         int_assert_o    
);

    // int
    localparam  S_INT_IDLE          = 4'b0001;
    localparam  S_INT_SYNC_ASSERT   = 4'b0010;
    localparam  S_INT_ASYNC_ASSERT  = 4'b0100;
    localparam  S_INT_MRET     = 4'b1000;

    // csr 
    localparam  S_CSR_IDLE          = 5'b00001;
    localparam  S_CSR_MSTATUS       = 5'b00010;
    localparam  S_CSR_MEPC          = 5'b00100;
    localparam  S_CSR_MSTATUS_MRET  = 5'b01000;
    localparam  S_CSR_MCAUSE        = 5'b10000;

    reg [3:0         ]           int_state;
    reg [4:0         ]           csr_state;
    reg [`InstAddrBus]           inst_addr;
    reg [31:0        ]           cause;


    assign hold_flag_o = ((int_state != S_INT_IDLE) | (csr_state != S_CSR_IDLE))? `HoldEnable: `HoldDisable;

    always @ (*) begin
        if (rst == `RstEnable ) begin
            int_state = S_INT_IDLE;
        end else begin
            if (inst_i == `INST_ECALL || inst_i == `INST_EBREAK ) begin
                if (div_started_i == `DivStop ) begin
                    int_state = S_INT_SYNC_ASSERT ;
                end else begin
                    int_state = S_INT_IDLE ;
                end
            end else if (int_flag_i != `INT_NONE && global_int_en_i == `True ) begin
                int_state = S_INT_ASYNC_ASSERT;
            end else if (inst_i == `INST_MRET ) begin
                int_state = S_INT_MRET;
            end else begin
                int_state = S_INT_IDLE;
            end
        end
    end


    always @ (posedge clk ) begin
        if (rst == `RstEnable) begin
            csr_state <= S_CSR_IDLE; 
            cause     <= `ZeroWord;
            inst_addr <= `ZeroWord;
        end else begin
            case (csr_state) 
                S_CSR_IDLE: begin
                    if (int_state == S_INT_SYNC_ASSERT) begin
                        csr_state <= S_CSR_MEPC;
                        if (jump_flag_i == `JumpEnable) begin
                            inst_addr <= jump_addr_i -4'h4;
                        end else begin
                            inst_addr <= inst_addr_i;
                        end
                        case (inst_i)
                            `INST_ECALL: begin
                                cause <= 32'd11;
                            end
                            `INST_EBREAK: begin
                                cause <= 32'd3;
                            end
                            default: begin
                                cause <= 32'd10;
                            end
                        endcase
                    end else if ( int_state == S_INT_ASYNC_ASSERT) begin
                        cause       <= 32'h80000004;
                        csr_state   <= S_CSR_MEPC;
                        if (jump_flag_i == `JumpEnable) begin
                            inst_addr <= jump_addr_i;
                        end else if (div_started_i == `DivStart) begin
                            inst_addr <= inst_addr_i -4'h4;
                        end else begin
                            inst_addr <= inst_addr_i;
                        end
                    end else if (int_state == S_INT_MRET) begin
                        csr_state <= S_CSR_MSTATUS_MRET;
                    end
                end
                S_CSR_MEPC: begin
                    csr_state <= S_CSR_MSTATUS;
                end
                S_CSR_MSTATUS: begin
                    csr_state <= S_CSR_MCAUSE;
                end
                S_CSR_MCAUSE: begin
                    csr_state <= S_CSR_IDLE;
                end
                S_CSR_MSTATUS_MRET: begin
                    csr_state <= S_CSR_IDLE;
                end
                default: begin
                    csr_state <= S_CSR_IDLE;   
                end
            endcase
        end
    end


    always @ (posedge clk) begin
        if (rst == `RstEnable) begin
            we_o    <= `WriteEnable;
            waddr_o <= `ZeroWord;
            data_o  <= `ZeroWord;
        end else begin
            case (csr_state)
                S_CSR_MEPC: begin
                    we_o    <= `WriteEnable;
                    waddr_o <= {20'h0, `CSR_MEPC};
                    data_o  <= inst_addr;
                end
                S_CSR_MCAUSE: begin
                    we_o    <= `WriteEnable;
                    waddr_o <= {20'h0, `CSR_MCAUSE};
                    data_o  <= cause;
                end
                S_CSR_MSTATUS: begin
                    we_o    <= `WriteEnable;
                    waddr_o <= {20'h0, `CSR_MSTATUS};
                    data_o  <= {csr_mstatus[31:4], 1'b0, csr_mstatus[2:0]};
                end
                S_CSR_MSTATUS_MRET: begin
                    we_o    <= `WriteEnable;
                    waddr_o <= {20'h0, `CSR_MSTATUS};
                    data_o  <= {csr_mstatus[31:4], csr_mstatus[7], csr_mstatus[2:0]};
                end
                default: begin
                    we_o    <= `WriteEnable;
                    waddr_o <= `ZeroWord;
                    data_o  <= `ZeroWord;
                end
            endcase
        end
    end

    always @ (posedge clk) begin
        if (rst == `RstEnable) begin
            int_assert_o    <= `INT_DEASSERT;
            int_addr_o      <= `ZeroWord;
        end else begin
            case (csr_state) 
                S_CSR_MCAUSE: begin
                     int_assert_o    <= `INT_ASSERT;                   
                     int_addr_o      <= csr_mtvec;
                end
                S_CSR_MSTATUS_MRET: begin
                     int_assert_o    <= `INT_ASSERT;                   
                     int_addr_o      <= csr_mepc;
                end
                default: begin
                    int_assert_o    <= `INT_DEASSERT;
                    int_addr_o      <= `ZeroWord;
                end
            endcase
        end
    end

endmodule
