`include "defines.v"
module ex (
    input   wire                rst,

    // from id
    input   wire    [`InstBus    ]  inst_i          ,
    input   wire    [`InstAddrBus]  inst_addr_i     ,
    input   wire                    reg_we_i        ,
    input   wire    [`RegAddrBus ]  reg_waddr_i     ,
    input   wire    [`RegBus     ]  reg1_rdata_i    ,
    input   wire    [`RegBus     ]  reg2_rdata_i    ,
    input   wire                    csr_we_i        ,
    input   wire    [`RegBus     ]  csr_rdata_i     ,
    input   wire    [`MemAddrBus ]  csr_waddr_i     ,
    input   wire                    int_assert_i    ,
    input   wire    [`InstAddrBus]  int_addr_i      ,
    input   wire    [`MemAddrBus ]  op1_i           ,
    input   wire    [`MemAddrBus ]  op2_i           ,
    input   wire    [`MemAddrBus ]  op1_jump_i      ,
    input   wire    [`MemAddrBus ]  op2_jump_i      ,

    // from mem
    input   wire    [`MemBus     ]  mem_rdata_i     ,

    // from div
    input   wire                    div_ready_i     ,
    input   wire    [`RegBus     ]  div_result_i    ,
    input   wire                    div_busy_i      ,
    input   wire    [`RegAddrBus ]  div_reg_waddr_i ,

    // to mem
    output  reg     [`MemBus     ]  mem_wdata_o     ,
    output  reg     [`MemAddrBus ]  mem_raddr_o     ,
    output  reg     [`MemAddrBus ]  mem_waddr_o     ,
    output  wire                    mem_we_o        ,
    output  wire                    mem_req_o       ,

    // to regs
    output  wire    [`RegBus     ]  reg_wdata_o     ,
    output  wire                    reg_we_o        ,
    output  wire    [`RegAddrBus ]  reg_waddr_o     ,
    
    // to csr reg
    output  reg     [`RegBus     ]  csr_wdata_o     ,
    output  wire                    csr_we_o        ,
    output  wire    [`MemAddrBus ]  csr_waddr_o     ,


    // to div
    output  wire                    div_start_o     ,
    output  reg     [`RegBus     ]  div_dividend_o  ,
    output  reg     [`RegBus     ]  div_divisor_o   ,   
    output  reg     [2:0         ]  div_op_o        ,
    output  reg     [`RegAddrBus ]  div_reg_waddr_o ,

    // to ctrl
    output  wire                    hold_flag_o     ,
    output  wire                    jump_flag_o     ,
    output  wire     [`InstAddrBus] jump_addr_o
    
    );
    wire    [1:0          ]  mem_raddr_index; 
    wire    [1:0          ]  mem_waddr_index; 
    wire    [`DoubleRegBus]  mul_temp; 
    wire    [`DoubleRegBus]  mul_temp_invert; 
    wire    [31:0         ]  sr_shift  ; 
    wire    [31:0         ]  sri_shift  ; 
    wire    [31:0         ]  sr_shift_mask  ; 
    wire    [31:0         ]  sri_shift_mask  ; 
    wire    [31:0         ]  op1_add_op2_res; 
    wire    [31:0         ]  op1_jump_add_op2_jump_res; 
    wire    [31:0         ]  reg1_data_invert  ; 
    wire    [31:0         ]  reg2_data_invert  ; 
    wire                     op1_ge_op2_signed;
    wire                     op1_ge_op2_unsigned;
    wire                     op1_eq_op2;
    reg     [`RegBus      ]  mul_op1;
    reg     [`RegBus      ]  mul_op2;
    wire    [6:0          ]  opcode; 
    wire    [2:0          ]  funct3; 
    wire    [6:0          ]  funct7; 
    wire    [4:0          ]  rd    ; 
    wire    [4:0          ]  uimm  ; 
    reg     [`RegBus      ]  reg_wdata;
    reg                      reg_we;
    reg     [`RegAddrBus  ]  reg_waddr;
    reg     [`RegBus      ]  div_wdata;
    reg                      div_we;
    reg     [`RegAddrBus  ]  div_waddr;
    reg                      div_hold_flag;
    reg                      div_jump_flag;
    reg     [`InstAddrBus]   div_jump_addr;
    reg                      hold_flag;
    reg                      jump_flag;
    reg     [`InstAddrBus]   jump_addr;
    reg                      mem_we;
    reg                      mem_req;
    reg                      div_start;


    assign  opcode = inst_i[6:0];
    assign  funct3 = inst_i[14:12];
    assign  funct7 = inst_i[31:25];
    assign  rd     = inst_i[11:7];
    assign  uimm   = inst_i[19:15];

    assign  sr_shift        = reg1_rdata_i  >> reg2_rdata_i[4:0];
    assign  sri_shift       = reg1_rdata_i  >> inst_i[24:20];
    assign  sr_shift_mask   = 32'hffffffff  >> reg2_rdata_i[4:0];
    assign  sri_shift_mask  = 32'hffffffff  >> inst_i[24:20];

    assign  op1_add_op2_res             = op1_i + op2_i;
    assign  op1_jump_add_op2_jump_res   = op1_jump_i + op2_jump_i;

    assign  reg1_data_invert = ~reg1_rdata_i + 1;
    assign  reg2_data_invert = ~reg2_rdata_i + 1;

    // comp
    assign  op1_ge_op2_signed   = $signed(op1_i) >= $signed(op2_i); 
    assign  op1_ge_op2_unsigned = op1_i >= op2_i; 
    assign  op1_eq_op2          = (op1_i == op2_i);

    assign  mul_temp        = mul_op1 * mul_op2;
    assign  mul_temp_invert = ~mul_temp + 1;

    assign  mem_raddr_index = (reg1_rdata_i + {{20{inst_i[31]}},inst_i[31:20]}) & 2'b11;
    assign  mem_waddr_index = (reg1_rdata_i + {{20{inst_i[31]}},inst_i[31:25], inst_i[11:7]}) & 2'b11;

    assign  div_start_o     = (int_assert_i == `INT_ASSERT)? `DivStop:div_start;

    assign  reg_wdata_o     = reg_wdata | div_wdata;


    assign  reg_we_o        = (int_assert_i == `INT_ASSERT)? `WriteDisable: (reg_we || div_we);
    assign  reg_waddr_o     = reg_waddr | div_waddr;

    assign  mem_we_o        = (int_assert_i == `INT_ASSERT)? `WriteDisable:mem_we;

    assign  mem_req_o       = (int_assert_i == `INT_ASSERT)? `RIB_NREQ:mem_req;






    assign  hold_flag_o     = hold_flag || div_hold_flag;
    assign  jump_flag_o     = jump_flag || div_jump_flag || ((int_assert_i == `INT_ASSERT)? `JumpEnable: `JumpDisable );
    assign  jump_addr_o     = (int_assert_i == `INT_ASSERT)? int_addr_i: (jump_addr | div_jump_addr);

    assign  csr_we_o        = (int_assert_i == `INT_ASSERT)? `WriteDisable: csr_we_i;
    assign  csr_waddr_o     = csr_waddr_i;




    // about mul inst
    always @ (*) begin
        if ((opcode == `INST_TYPE_R_M) && (funct7 == 7'b0000001)) begin
            case (funct3)
                `INST_MUL,`INST_MULHU: begin
                    mul_op1 = reg1_rdata_i;
                    mul_op2 = reg2_rdata_i;
                end
                `INST_MULHSU: begin
                    mul_op1 = (reg1_rdata_i[31] == 1'b1)? (reg1_data_invert):reg1_rdata_i;
                    mul_op2 = reg2_rdata_i;
                end
                `INST_MULH: begin
                    mul_op1 = (reg1_rdata_i[31] == 1'b1)? (reg1_data_invert):reg1_rdata_i;
                    mul_op2 = (reg2_rdata_i[31] == 2'b1)? (reg2_data_invert):reg2_rdata_i;
                end
                default: begin
                    mul_op1 = reg1_rdata_i;
                    mul_op2 = reg2_rdata_i;
                end
            endcase
        end else begin
            mul_op1 = reg1_rdata_i;
            mul_op2 = reg2_rdata_i;
        end
    end

    // about div inst
    always @ (*)begin
        div_dividend_o = reg1_rdata_i;
        div_divisor_o  = reg2_rdata_i;
        div_op_o       = funct3;
        div_reg_waddr_o= reg_waddr_i;
        if ((opcode == `INST_TYPE_R_M) && (funct7 == 7'b0000001)) begin
            div_we      = `WriteDisable;
            div_wdata   = `ZeroWord  ;
            div_waddr   = `ZeroWord  ;
            case (funct3)
                `INST_DIV, `INST_DIVU, `INST_REM, `INST_REMU: begin
                    div_start       = `DivStart;
                    div_jump_flag   = `JumpEnable ;
                    div_hold_flag   = `HoldEnable;
                    div_jump_addr   = op1_jump_add_op2_jump_res;
                end
                default: begin
                    div_start       = `DivStop ;
                    div_jump_flag   = `JumpDisable;
                    div_hold_flag   = `HoldDisable;
                    div_jump_addr   = `ZeroWord;
                end
            endcase
        end else begin
            div_jump_flag   = `JumpDisable;
            div_jump_addr   = `ZeroWord;
            if (div_busy_i == `True ) begin
                div_start       = `DivStart;
                div_we          = `WriteDisable;
                div_wdata       = `ZeroWord  ;
                div_waddr       = `ZeroWord  ;
                div_hold_flag   = `HoldEnable;
            end else begin
                div_start       = `DivStop ;
                div_hold_flag   = `HoldDisable;
                if (div_ready_i == `DivResultReady) begin
                    div_we          = `WriteEnable;
                    div_wdata       = div_result_i;
                    div_waddr       = div_reg_waddr_i  ;
                end else begin
                    div_we          = `WriteDisable;
                    div_wdata       = `ZeroWord  ;
                    div_waddr       = `ZeroWord  ;
                end
            end
        end
    end

    // ex
    always @ (*) begin
        reg_we      = reg_we_i;
        reg_waddr   = reg_waddr_i;
        mem_req     = `RIB_NREQ ;
        csr_wdata_o = `ZeroWord ;
        
        case (opcode)
            `INST_TYPE_I: begin
                case (funct3) 
                    `INST_ADDI: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = op1_add_op2_res;
                    end
                    `INST_SLTI: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = {32{(~op1_ge_op2_signed)}} & 32'h1;
                    end
                    `INST_SLTIU: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = {32{(~op1_ge_op2_unsigned)}} & 32'h1;
                    end
                    `INST_XORI: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = op1_i ^ op2_i;
                    end
                    `INST_ORI: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = op1_i | op2_i;
                    end
                    `INST_ANDI: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = op1_i & op2_i;
                    end
                    `INST_SLLI: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = reg1_rdata_i << inst_i[24:20];
                    end
                    `INST_SRI: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        if (inst_i[30] == 1'b1) begin
                            reg_wdata   = (sri_shift & sri_shift_mask) | ({32{reg1_rdata_i[31]}} & (~sri_shift_mask));
                        end else begin
                            reg_wdata   = reg1_rdata_i >> inst_i[24:20];
                        end 
                    end
                    default: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = `ZeroWord  ;
                    end
                endcase
            end
            `INST_TYPE_R_M: begin
                if ((funct7 == 7'b0000000) || (funct7 == 7'b0100000)) begin
                    case (funct3)
                        `INST_ADD_SUB: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            if (inst_i[30] == 1'b0) begin
                                reg_wdata   = op1_add_op2_res  ;
                            end else begin
                                reg_wdata   = op1_i-op2_i  ;
                            end
                        end
                        `INST_SLL: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = op1_i << op2_i[4:0];
                        end
                        `INST_SLT: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = {32{(~op1_ge_op2_signed)}} & 32'h1;
                        end
                        `INST_SLTU: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = {32{(~op1_ge_op2_unsigned)}} & 32'h1;
                        end
                        `INST_XOR: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = op1_i ^ op2_i;
                        end
                        `INST_SR: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            if (inst_i[30] == 1'b1) begin
                                reg_wdata   = (sr_shift & sr_shift_mask) | ({32{reg1_rdata_i[31]}} & (~sr_shift_mask));
                            end else begin
                                 reg_wdata   = reg1_rdata_i >> reg2_rdata_i[4:0];                                                    
                            end
                        end
                        `INST_OR: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = op1_i | op2_i;
                        end
                        `INST_AND: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = op1_i & op2_i;
                        end
                        default: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = `ZeroWord  ;
                        end
                    endcase
                end else if(funct7 == 7'b0000001) begin
                    case (funct3)
                        `INST_MUL   : begin 
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = mul_temp[31:0];
                        end
                        `INST_MULHU : begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = mul_temp[63:32];
                        end
                        `INST_MULH: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            case ({reg1_rdata_i[31], reg2_rdata_i[31]}) 
                                2'b00: begin
                                    reg_wdata   = mul_temp[63:32];
                                end
                                2'b11: begin
                                    reg_wdata   = mul_temp[63:32];
                                end
                                2'b10: begin
                                    reg_wdata   = mul_temp_invert[63:32];
                                end
                                default: begin
                                    reg_wdata   = mul_temp_invert[63:32];
                                end
                            endcase
                        end
                        `INST_MULHSU : begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            if (reg1_rdata_i[31] == 1'b1) begin
                                reg_wdata   = mul_temp_invert[63:32];
                            end else begin
                                reg_wdata   = mul_temp[63:32];
                            end
                        end
                        default: begin
                            jump_flag   = `JumpDisable;
                            hold_flag   = `HoldDisable;
                            jump_addr   = `ZeroWord  ;
                            mem_wdata_o = `ZeroWord  ;
                            mem_raddr_o = `ZeroWord  ;     
                            mem_waddr_o = `ZeroWord  ;     
                            mem_we      = `WriteDisable;
                            reg_wdata   = `ZeroWord  ;
                        end
                    endcase
                end else begin
                    jump_flag   = `JumpDisable;
                    hold_flag   = `HoldDisable;
                    jump_addr   = `ZeroWord  ;
                    mem_wdata_o = `ZeroWord  ;
                    mem_raddr_o = `ZeroWord  ;     
                    mem_waddr_o = `ZeroWord  ;     
                    mem_we      = `WriteDisable;
                    reg_wdata   = `ZeroWord  ;
                end
            end
            `INST_TYPE_L: begin
                case (funct3)
                    `INST_LB : begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        mem_req     = `RIB_REQ;
                        mem_raddr_o = op1_add_op2_res;
                        case (mem_raddr_index)
                            2'b00: begin
                                reg_wdata   = {{24{mem_rdata_i[7]}}, mem_rdata_i[7:0]};
                            end
                            2'b01: begin
                                reg_wdata   = {{24{mem_rdata_i[15]}}, mem_rdata_i[15:8]};
                            end
                            2'b10: begin
                                reg_wdata   = {{24{mem_rdata_i[23]}}, mem_rdata_i[23:16]};
                            end
                            default: begin
                                reg_wdata   = {{24{mem_rdata_i[31]}}, mem_rdata_i[31:24]};
                            end
                        endcase
                    end
                    `INST_LH : begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        mem_req     = `RIB_REQ;
                        mem_raddr_o = op1_add_op2_res;
                        if (mem_raddr_index == 2'b0) begin
                            reg_wdata   = {{16{mem_rdata_i[15]}}, mem_rdata_i[15:0]};
                        end else begin
                            reg_wdata   = {{16{mem_rdata_i[31]}}, mem_rdata_i[31:16]};
                        end
                    end
                    `INST_LW : begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        mem_req     = `RIB_REQ;
                        mem_raddr_o = op1_add_op2_res;
                        reg_wdata   = mem_rdata_i;
                    end
                    `INST_LBU : begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        mem_req     = `RIB_REQ;
                        mem_raddr_o = op1_add_op2_res;
                        case (mem_raddr_index)
                            2'b00: begin
                                reg_wdata   = {24'h0, mem_rdata_i[7:0]};
                            end
                            2'b01: begin
                                reg_wdata   = {24'h0, mem_rdata_i[15:8]};
                            end
                            2'b10: begin
                                reg_wdata   = {24'h0, mem_rdata_i[23:16]};
                            end
                            default: begin
                                reg_wdata   = {24'h0, mem_rdata_i[31:24]};
                            end
                        endcase
                    end
                    `INST_LHU : begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        mem_req     = `RIB_REQ;
                        mem_raddr_o = op1_add_op2_res;
                        if (mem_raddr_index == 2'b0) begin
                            reg_wdata   = {16'h0, mem_rdata_i[15:0]};
                        end else begin
                            reg_wdata   = {16'h0, mem_rdata_i[31:16]};
                        end
                    end
                    default: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = `ZeroWord  ;
                    end
                endcase
            end
            `INST_TYPE_S: begin
                case (funct3)
                    `INST_SB: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable; 
                        jump_addr   = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        mem_we      = `WriteEnable;
                        mem_req     = `RIB_REQ;
                        mem_wdata_o = op1_add_op2_res  ;
                        mem_raddr_o = op1_add_op2_res  ;    
                        case (mem_waddr_index)
                            2'b00: begin
                                mem_waddr_o = {mem_rdata_i[31:8], reg2_rdata_i[7:0]};
                            end
                            2'b01: begin
                                mem_waddr_o = {mem_rdata_i[31:16], reg2_rdata_i[7:0], mem_rdata_i[7:0]};
                            end
                            2'b10: begin
                                mem_waddr_o = {mem_rdata_i[31:24], reg2_rdata_i[7:0], mem_rdata_i[15:0]};
                            end
                            default: begin
                                mem_waddr_o = {reg2_rdata_i[7:0], mem_rdata_i[23:0]};
                            end
                        endcase
                    end
                    `INST_SH: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable; 
                        jump_addr   = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        mem_we      = `WriteEnable;
                        mem_req     = `RIB_REQ;
                        mem_wdata_o = op1_add_op2_res  ;
                        mem_raddr_o = op1_add_op2_res  ;
                        if (mem_waddr_index == 2'b00) begin
                            mem_waddr_o = {mem_rdata_i[31:16], reg2_rdata_i[15:0]};
                        end else begin
                            mem_waddr_o = {reg2_rdata_i[15:0], mem_rdata_i[15:0]};
                        end
                    end
                    `INST_SW: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable; 
                        jump_addr   = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        mem_we      = `WriteEnable;                         
                        mem_req     = `RIB_REQ;
                        mem_wdata_o = op1_add_op2_res  ;
                        mem_raddr_o = op1_add_op2_res  ;
                        mem_waddr_o = reg2_rdata_i;
                    end
                    default : begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable; 
                        jump_addr   = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        mem_we      = `WriteDisable;                         
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;
                    end
                endcase
            end
            `INST_TYPE_B: begin
                case (funct3)
                    `INST_BEQ : begin
                        hold_flag   = `HoldDisable; 
                        mem_we      = `WriteDisable;                         
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        jump_flag   = op1_eq_op2 & `JumpEnable; 
                        jump_addr   = {32{op1_eq_op2}} & op1_jump_add_op2_jump_res;
                    end
                    `INST_BNE : begin
                        hold_flag   = `HoldDisable; 
                        mem_we      = `WriteDisable;                         
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        jump_flag   = (~op1_eq_op2) & `JumpEnable; 
                        jump_addr   = {32{(~op1_eq_op2)}} & op1_jump_add_op2_jump_res;
                    end
                    `INST_BLT : begin
                        hold_flag   = `HoldDisable; 
                        mem_we      = `WriteDisable;                         
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        jump_flag   = (~op1_ge_op2_signed) & `JumpEnable; 
                        jump_addr   = {32{(~op1_ge_op2_signed)}} & op1_jump_add_op2_jump_res;
                    end
                    `INST_BGE : begin
                        hold_flag   = `HoldDisable; 
                        mem_we      = `WriteDisable;                         
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        jump_flag   = (op1_ge_op2_signed) & `JumpEnable; 
                        jump_addr   = {32{(op1_ge_op2_signed)}} & op1_jump_add_op2_jump_res;
                    end
                    `INST_BLTU: begin
                        hold_flag   = `HoldDisable; 
                        mem_we      = `WriteDisable;                         
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        jump_flag   = (~op1_ge_op2_unsigned) & `JumpEnable; 
                        jump_addr   = {32{(~op1_ge_op2_unsigned)}} & op1_jump_add_op2_jump_res;
                    end
                    `INST_BGEU: begin 
                        hold_flag   = `HoldDisable; 
                        mem_we      = `WriteDisable;                         
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;
                        mem_waddr_o = `ZeroWord  ;
                        reg_wdata   = `ZeroWord  ;
                        jump_flag   = (op1_ge_op2_unsigned) & `JumpEnable; 
                        jump_addr   = {32{(op1_ge_op2_unsigned)}} & op1_jump_add_op2_jump_res;
                    end
                    default: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = `ZeroWord  ;
                    end
                endcase
            end
            `INST_JAL, `INST_JALR: begin
                jump_flag   = `JumpEnable;
                hold_flag   = `HoldDisable;
                jump_addr   = op1_jump_add_op2_jump_res  ;
                mem_wdata_o = `ZeroWord  ;
                mem_raddr_o = `ZeroWord  ;     
                mem_waddr_o = `ZeroWord  ;     
                mem_we      = `WriteDisable;
                reg_wdata   = op1_add_op2_res  ;
            end
            `INST_LUI, `INST_AUIPC: begin
                jump_flag   = `JumpDisable;
                hold_flag   = `HoldDisable;
                jump_addr   = `ZeroWord  ;
                mem_wdata_o = `ZeroWord  ;
                mem_raddr_o = `ZeroWord  ;     
                mem_waddr_o = `ZeroWord  ;     
                mem_we      = `WriteDisable;
                reg_wdata   = op1_add_op2_res  ;
            end
            `INST_NOP_OP: begin
                jump_flag   = `JumpDisable;
                hold_flag   = `HoldDisable;
                jump_addr   = `ZeroWord  ;
                mem_wdata_o = `ZeroWord  ;
                mem_raddr_o = `ZeroWord  ;     
                mem_waddr_o = `ZeroWord  ;     
                mem_we      = `WriteDisable;
                reg_wdata   = `ZeroWord  ;
            end
            `INST_FENCE: begin
                jump_flag   = `JumpEnable;
                hold_flag   = `HoldDisable;
                jump_addr   = op1_jump_add_op2_jump_res  ;
                mem_wdata_o = `ZeroWord  ;
                mem_raddr_o = `ZeroWord  ;     
                mem_waddr_o = `ZeroWord  ;     
                mem_we      = `WriteDisable;
                reg_wdata   = `ZeroWord  ;
            end
            `INST_CSR: begin
                jump_flag   = `JumpDisable;
                hold_flag   = `HoldDisable;
                jump_addr   = `ZeroWord  ;
                mem_wdata_o = `ZeroWord  ;
                mem_raddr_o = `ZeroWord  ;     
                mem_waddr_o = `ZeroWord  ;     
                mem_we      = `WriteDisable;
                case (funct3)
                    `INST_CSRRW : begin
                        csr_wdata_o = reg1_rdata_i;
                        reg_wdata   = csr_rdata_i;
                    end
                    `INST_CSRRS : begin
                        csr_wdata_o = reg1_rdata_i | csr_rdata_i;
                        reg_wdata   = csr_rdata_i;
                    end
                    `INST_CSRRC : begin
                        csr_wdata_o = (~reg1_rdata_i) | csr_rdata_i;
                        reg_wdata   = csr_rdata_i;
                    end
                    `INST_CSRRWI: begin
                        csr_wdata_o = {27'h0, uimm};
                        reg_wdata   = csr_rdata_i;
                    end
                    `INST_CSRRSI: begin
                        csr_wdata_o = {27'h0, uimm} | csr_rdata_i;
                        reg_wdata   = csr_rdata_i;
                    end
                    `INST_CSRRCI:begin
                        csr_wdata_o = (~{27'h0, uimm}) & csr_rdata_i;
                        reg_wdata   = csr_rdata_i;
                    end
                    default: begin
                        jump_flag   = `JumpDisable;
                        hold_flag   = `HoldDisable;
                        jump_addr   = `ZeroWord  ;
                        mem_wdata_o = `ZeroWord  ;
                        mem_raddr_o = `ZeroWord  ;     
                        mem_waddr_o = `ZeroWord  ;     
                        mem_we      = `WriteDisable;
                        reg_wdata   = `ZeroWord  ;
                    end
                endcase
            end
            default: begin
                jump_flag   = `JumpDisable;
                hold_flag   = `HoldDisable;
                jump_addr   = `ZeroWord  ;
                mem_wdata_o = `ZeroWord  ;
                mem_raddr_o = `ZeroWord  ;     
                mem_waddr_o = `ZeroWord  ;     
                mem_we      = `WriteDisable;
                reg_wdata   = `ZeroWord  ;
            end
        endcase
    end


endmodule
